`include "src/float/div.v"

module tb();

wire [31:0] s;
reg [31:0] a, b;
wire ze;

divf df(s, ze, a, b);

initial begin
$monitor("%b %b %b %b\n", df.ssign, df.sexp, df.smant, s);
//3.2. -1.3
a = 32'b01000000010011001100110011001101;
b = 32'b10111111101001100110011001100110;
#100;
$display("11000000000111011000100111011001");
//1, 5
a = 32'b00111111100000000000000000000000;
b = 32'b01000000101000000000000000000000;
#100;
$display("00111110010011001100110011001101");
//-5, 3
a = 32'b11000000101000000000000000000000;
b = 32'b01000000010000000000000000000000;
#100;
$display("10111111110101010101010101010101");
//-3, -3.6
a = 32'b11000000010000000000000000000000;
b = 32'b11000000011001100110011001100110;
#100;
$display("00111111010101010101010101010101");
//4.153844e34, 4.153844e34
a = 32'b01111001000000000000000000001101;
b = 32'b01111001000000000000000000001101;
#100;
$display("00111111100000000000000000000000");
end

endmodule