`include "src/float/add.v"

module tb();

wire [31:0] s;
reg [31:0] a, b;

addf af(s, a, b);

initial begin
$monitor("%b %b %b %b\n", af.aexp, af.bexp, af.smant, s);
//3.2. -1.3
a = 32'b01000000010011001100110011001101;
b = 32'b10111111101001100110011001100110;
#100;
$display("00111111111100110011001100110011");
//3.2. 1.3
a = 32'b01000000010011001100110011001101;
b = 32'b00111111101001100110011001100110;
#100;
$display("01000000100100000000000000000000");
//1, 5
a = 32'b00111111100000000000000000000000;
b = 32'b01000000101000000000000000000000;
#100;
$display("01000000110000000000000000000000");
//69, 5
a = 32'b01000010100010100000000000000000;
b = 32'b01000000101000000000000000000000;
#100;
$display("01000010100101000000000000000000");
//2.3, -2.3
a = 32'b01000000000100110011001100110011;
b = 32'b11000000000100110011001100110011;
#100;
$display("0");
//5, -2.3
a = 32'b01000000101000000000000000000000;
b = 32'b11000000000100110011001100110011;
#100;
$display("01000000001011001100110011001101");
$finish;
end

endmodule
